module forwarding_unit(input ex_control_i,
							  input wb_control_i,
							  output[1:0] rs_muxcontrol_o,
							  output[1:0] rt_muxcontrol_o);
							  
							  
endmodule