module pipelineEMWB(input in_i,
								output out_o);
								
								
								
								
endmodule